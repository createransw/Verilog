module mux64_4_2(y0, y1, y2, y3, x, z);

    input wire[63:0] y0;
    input wire[63:0] y1;
    input wire[63:0] y2;
    input wire[63:0] y3;

    input wire[1:0] x;

    output wire[63:0] z;

    wire[1:0] inv;
    not i0(inv[0], x[0]);
    not i1(inv[1], x[1]);

    wire[63 : 0] first_0;
    wire[63 : 0] first_1;

    and f_00(first_0[0], y0[0], inv[0]);
    and f_10(first_1[0], y1[0], x[0]);
    and f_01(first_0[1], y0[1], inv[0]);
    and f_11(first_1[1], y1[1], x[0]);
    and f_02(first_0[2], y0[2], inv[0]);
    and f_12(first_1[2], y1[2], x[0]);
    and f_03(first_0[3], y0[3], inv[0]);
    and f_13(first_1[3], y1[3], x[0]);
    and f_04(first_0[4], y0[4], inv[0]);
    and f_14(first_1[4], y1[4], x[0]);
    and f_05(first_0[5], y0[5], inv[0]);
    and f_15(first_1[5], y1[5], x[0]);
    and f_06(first_0[6], y0[6], inv[0]);
    and f_16(first_1[6], y1[6], x[0]);
    and f_07(first_0[7], y0[7], inv[0]);
    and f_17(first_1[7], y1[7], x[0]);
    and f_08(first_0[8], y0[8], inv[0]);
    and f_18(first_1[8], y1[8], x[0]);
    and f_09(first_0[9], y0[9], inv[0]);
    and f_19(first_1[9], y1[9], x[0]);
    and f_010(first_0[10], y0[10], inv[0]);
    and f_110(first_1[10], y1[10], x[0]);
    and f_011(first_0[11], y0[11], inv[0]);
    and f_111(first_1[11], y1[11], x[0]);
    and f_012(first_0[12], y0[12], inv[0]);
    and f_112(first_1[12], y1[12], x[0]);
    and f_013(first_0[13], y0[13], inv[0]);
    and f_113(first_1[13], y1[13], x[0]);
    and f_014(first_0[14], y0[14], inv[0]);
    and f_114(first_1[14], y1[14], x[0]);
    and f_015(first_0[15], y0[15], inv[0]);
    and f_115(first_1[15], y1[15], x[0]);
    and f_016(first_0[16], y0[16], inv[0]);
    and f_116(first_1[16], y1[16], x[0]);
    and f_017(first_0[17], y0[17], inv[0]);
    and f_117(first_1[17], y1[17], x[0]);
    and f_018(first_0[18], y0[18], inv[0]);
    and f_118(first_1[18], y1[18], x[0]);
    and f_019(first_0[19], y0[19], inv[0]);
    and f_119(first_1[19], y1[19], x[0]);
    and f_020(first_0[20], y0[20], inv[0]);
    and f_120(first_1[20], y1[20], x[0]);
    and f_021(first_0[21], y0[21], inv[0]);
    and f_121(first_1[21], y1[21], x[0]);
    and f_022(first_0[22], y0[22], inv[0]);
    and f_122(first_1[22], y1[22], x[0]);
    and f_023(first_0[23], y0[23], inv[0]);
    and f_123(first_1[23], y1[23], x[0]);
    and f_024(first_0[24], y0[24], inv[0]);
    and f_124(first_1[24], y1[24], x[0]);
    and f_025(first_0[25], y0[25], inv[0]);
    and f_125(first_1[25], y1[25], x[0]);
    and f_026(first_0[26], y0[26], inv[0]);
    and f_126(first_1[26], y1[26], x[0]);
    and f_027(first_0[27], y0[27], inv[0]);
    and f_127(first_1[27], y1[27], x[0]);
    and f_028(first_0[28], y0[28], inv[0]);
    and f_128(first_1[28], y1[28], x[0]);
    and f_029(first_0[29], y0[29], inv[0]);
    and f_129(first_1[29], y1[29], x[0]);
    and f_030(first_0[30], y0[30], inv[0]);
    and f_130(first_1[30], y1[30], x[0]);
    and f_031(first_0[31], y0[31], inv[0]);
    and f_131(first_1[31], y1[31], x[0]);
    and f_032(first_0[32], y0[32], inv[0]);
    and f_132(first_1[32], y1[32], x[0]);
    and f_033(first_0[33], y0[33], inv[0]);
    and f_133(first_1[33], y1[33], x[0]);
    and f_034(first_0[34], y0[34], inv[0]);
    and f_134(first_1[34], y1[34], x[0]);
    and f_035(first_0[35], y0[35], inv[0]);
    and f_135(first_1[35], y1[35], x[0]);
    and f_036(first_0[36], y0[36], inv[0]);
    and f_136(first_1[36], y1[36], x[0]);
    and f_037(first_0[37], y0[37], inv[0]);
    and f_137(first_1[37], y1[37], x[0]);
    and f_038(first_0[38], y0[38], inv[0]);
    and f_138(first_1[38], y1[38], x[0]);
    and f_039(first_0[39], y0[39], inv[0]);
    and f_139(first_1[39], y1[39], x[0]);
    and f_040(first_0[40], y0[40], inv[0]);
    and f_140(first_1[40], y1[40], x[0]);
    and f_041(first_0[41], y0[41], inv[0]);
    and f_141(first_1[41], y1[41], x[0]);
    and f_042(first_0[42], y0[42], inv[0]);
    and f_142(first_1[42], y1[42], x[0]);
    and f_043(first_0[43], y0[43], inv[0]);
    and f_143(first_1[43], y1[43], x[0]);
    and f_044(first_0[44], y0[44], inv[0]);
    and f_144(first_1[44], y1[44], x[0]);
    and f_045(first_0[45], y0[45], inv[0]);
    and f_145(first_1[45], y1[45], x[0]);
    and f_046(first_0[46], y0[46], inv[0]);
    and f_146(first_1[46], y1[46], x[0]);
    and f_047(first_0[47], y0[47], inv[0]);
    and f_147(first_1[47], y1[47], x[0]);
    and f_048(first_0[48], y0[48], inv[0]);
    and f_148(first_1[48], y1[48], x[0]);
    and f_049(first_0[49], y0[49], inv[0]);
    and f_149(first_1[49], y1[49], x[0]);
    and f_050(first_0[50], y0[50], inv[0]);
    and f_150(first_1[50], y1[50], x[0]);
    and f_051(first_0[51], y0[51], inv[0]);
    and f_151(first_1[51], y1[51], x[0]);
    and f_052(first_0[52], y0[52], inv[0]);
    and f_152(first_1[52], y1[52], x[0]);
    and f_053(first_0[53], y0[53], inv[0]);
    and f_153(first_1[53], y1[53], x[0]);
    and f_054(first_0[54], y0[54], inv[0]);
    and f_154(first_1[54], y1[54], x[0]);
    and f_055(first_0[55], y0[55], inv[0]);
    and f_155(first_1[55], y1[55], x[0]);
    and f_056(first_0[56], y0[56], inv[0]);
    and f_156(first_1[56], y1[56], x[0]);
    and f_057(first_0[57], y0[57], inv[0]);
    and f_157(first_1[57], y1[57], x[0]);
    and f_058(first_0[58], y0[58], inv[0]);
    and f_158(first_1[58], y1[58], x[0]);
    and f_059(first_0[59], y0[59], inv[0]);
    and f_159(first_1[59], y1[59], x[0]);
    and f_060(first_0[60], y0[60], inv[0]);
    and f_160(first_1[60], y1[60], x[0]);
    and f_061(first_0[61], y0[61], inv[0]);
    and f_161(first_1[61], y1[61], x[0]);
    and f_062(first_0[62], y0[62], inv[0]);
    and f_162(first_1[62], y1[62], x[0]);
    and f_063(first_0[63], y0[63], inv[0]);
    and f_163(first_1[63], y1[63], x[0]);

    wire[63 : 0] first;

    or f0(first[0], first_0[0], first_1[0]);
    or f1(first[1], first_0[1], first_1[1]);
    or f2(first[2], first_0[2], first_1[2]);
    or f3(first[3], first_0[3], first_1[3]);
    or f4(first[4], first_0[4], first_1[4]);
    or f5(first[5], first_0[5], first_1[5]);
    or f6(first[6], first_0[6], first_1[6]);
    or f7(first[7], first_0[7], first_1[7]);
    or f8(first[8], first_0[8], first_1[8]);
    or f9(first[9], first_0[9], first_1[9]);
    or f10(first[10], first_0[10], first_1[10]);
    or f11(first[11], first_0[11], first_1[11]);
    or f12(first[12], first_0[12], first_1[12]);
    or f13(first[13], first_0[13], first_1[13]);
    or f14(first[14], first_0[14], first_1[14]);
    or f15(first[15], first_0[15], first_1[15]);
    or f16(first[16], first_0[16], first_1[16]);
    or f17(first[17], first_0[17], first_1[17]);
    or f18(first[18], first_0[18], first_1[18]);
    or f19(first[19], first_0[19], first_1[19]);
    or f20(first[20], first_0[20], first_1[20]);
    or f21(first[21], first_0[21], first_1[21]);
    or f22(first[22], first_0[22], first_1[22]);
    or f23(first[23], first_0[23], first_1[23]);
    or f24(first[24], first_0[24], first_1[24]);
    or f25(first[25], first_0[25], first_1[25]);
    or f26(first[26], first_0[26], first_1[26]);
    or f27(first[27], first_0[27], first_1[27]);
    or f28(first[28], first_0[28], first_1[28]);
    or f29(first[29], first_0[29], first_1[29]);
    or f30(first[30], first_0[30], first_1[30]);
    or f31(first[31], first_0[31], first_1[31]);
    or f32(first[32], first_0[32], first_1[32]);
    or f33(first[33], first_0[33], first_1[33]);
    or f34(first[34], first_0[34], first_1[34]);
    or f35(first[35], first_0[35], first_1[35]);
    or f36(first[36], first_0[36], first_1[36]);
    or f37(first[37], first_0[37], first_1[37]);
    or f38(first[38], first_0[38], first_1[38]);
    or f39(first[39], first_0[39], first_1[39]);
    or f40(first[40], first_0[40], first_1[40]);
    or f41(first[41], first_0[41], first_1[41]);
    or f42(first[42], first_0[42], first_1[42]);
    or f43(first[43], first_0[43], first_1[43]);
    or f44(first[44], first_0[44], first_1[44]);
    or f45(first[45], first_0[45], first_1[45]);
    or f46(first[46], first_0[46], first_1[46]);
    or f47(first[47], first_0[47], first_1[47]);
    or f48(first[48], first_0[48], first_1[48]);
    or f49(first[49], first_0[49], first_1[49]);
    or f50(first[50], first_0[50], first_1[50]);
    or f51(first[51], first_0[51], first_1[51]);
    or f52(first[52], first_0[52], first_1[52]);
    or f53(first[53], first_0[53], first_1[53]);
    or f54(first[54], first_0[54], first_1[54]);
    or f55(first[55], first_0[55], first_1[55]);
    or f56(first[56], first_0[56], first_1[56]);
    or f57(first[57], first_0[57], first_1[57]);
    or f58(first[58], first_0[58], first_1[58]);
    or f59(first[59], first_0[59], first_1[59]);
    or f60(first[60], first_0[60], first_1[60]);
    or f61(first[61], first_0[61], first_1[61]);
    or f62(first[62], first_0[62], first_1[62]);
    or f63(first[63], first_0[63], first_1[63]);

    wire[63 : 0] second_0;
    wire[63 : 0] second_1;

    and s_00(second_0[0], y2[0], inv[0]);
    and s_10(second_1[0], y3[0], x[0]);
    and s_01(second_0[1], y2[1], inv[0]);
    and s_11(second_1[1], y3[1], x[0]);
    and s_02(second_0[2], y2[2], inv[0]);
    and s_12(second_1[2], y3[2], x[0]);
    and s_03(second_0[3], y2[3], inv[0]);
    and s_13(second_1[3], y3[3], x[0]);
    and s_04(second_0[4], y2[4], inv[0]);
    and s_14(second_1[4], y3[4], x[0]);
    and s_05(second_0[5], y2[5], inv[0]);
    and s_15(second_1[5], y3[5], x[0]);
    and s_06(second_0[6], y2[6], inv[0]);
    and s_16(second_1[6], y3[6], x[0]);
    and s_07(second_0[7], y2[7], inv[0]);
    and s_17(second_1[7], y3[7], x[0]);
    and s_08(second_0[8], y2[8], inv[0]);
    and s_18(second_1[8], y3[8], x[0]);
    and s_09(second_0[9], y2[9], inv[0]);
    and s_19(second_1[9], y3[9], x[0]);
    and s_010(second_0[10], y2[10], inv[0]);
    and s_110(second_1[10], y3[10], x[0]);
    and s_011(second_0[11], y2[11], inv[0]);
    and s_111(second_1[11], y3[11], x[0]);
    and s_012(second_0[12], y2[12], inv[0]);
    and s_112(second_1[12], y3[12], x[0]);
    and s_013(second_0[13], y2[13], inv[0]);
    and s_113(second_1[13], y3[13], x[0]);
    and s_014(second_0[14], y2[14], inv[0]);
    and s_114(second_1[14], y3[14], x[0]);
    and s_015(second_0[15], y2[15], inv[0]);
    and s_115(second_1[15], y3[15], x[0]);
    and s_016(second_0[16], y2[16], inv[0]);
    and s_116(second_1[16], y3[16], x[0]);
    and s_017(second_0[17], y2[17], inv[0]);
    and s_117(second_1[17], y3[17], x[0]);
    and s_018(second_0[18], y2[18], inv[0]);
    and s_118(second_1[18], y3[18], x[0]);
    and s_019(second_0[19], y2[19], inv[0]);
    and s_119(second_1[19], y3[19], x[0]);
    and s_020(second_0[20], y2[20], inv[0]);
    and s_120(second_1[20], y3[20], x[0]);
    and s_021(second_0[21], y2[21], inv[0]);
    and s_121(second_1[21], y3[21], x[0]);
    and s_022(second_0[22], y2[22], inv[0]);
    and s_122(second_1[22], y3[22], x[0]);
    and s_023(second_0[23], y2[23], inv[0]);
    and s_123(second_1[23], y3[23], x[0]);
    and s_024(second_0[24], y2[24], inv[0]);
    and s_124(second_1[24], y3[24], x[0]);
    and s_025(second_0[25], y2[25], inv[0]);
    and s_125(second_1[25], y3[25], x[0]);
    and s_026(second_0[26], y2[26], inv[0]);
    and s_126(second_1[26], y3[26], x[0]);
    and s_027(second_0[27], y2[27], inv[0]);
    and s_127(second_1[27], y3[27], x[0]);
    and s_028(second_0[28], y2[28], inv[0]);
    and s_128(second_1[28], y3[28], x[0]);
    and s_029(second_0[29], y2[29], inv[0]);
    and s_129(second_1[29], y3[29], x[0]);
    and s_030(second_0[30], y2[30], inv[0]);
    and s_130(second_1[30], y3[30], x[0]);
    and s_031(second_0[31], y2[31], inv[0]);
    and s_131(second_1[31], y3[31], x[0]);
    and s_032(second_0[32], y2[32], inv[0]);
    and s_132(second_1[32], y3[32], x[0]);
    and s_033(second_0[33], y2[33], inv[0]);
    and s_133(second_1[33], y3[33], x[0]);
    and s_034(second_0[34], y2[34], inv[0]);
    and s_134(second_1[34], y3[34], x[0]);
    and s_035(second_0[35], y2[35], inv[0]);
    and s_135(second_1[35], y3[35], x[0]);
    and s_036(second_0[36], y2[36], inv[0]);
    and s_136(second_1[36], y3[36], x[0]);
    and s_037(second_0[37], y2[37], inv[0]);
    and s_137(second_1[37], y3[37], x[0]);
    and s_038(second_0[38], y2[38], inv[0]);
    and s_138(second_1[38], y3[38], x[0]);
    and s_039(second_0[39], y2[39], inv[0]);
    and s_139(second_1[39], y3[39], x[0]);
    and s_040(second_0[40], y2[40], inv[0]);
    and s_140(second_1[40], y3[40], x[0]);
    and s_041(second_0[41], y2[41], inv[0]);
    and s_141(second_1[41], y3[41], x[0]);
    and s_042(second_0[42], y2[42], inv[0]);
    and s_142(second_1[42], y3[42], x[0]);
    and s_043(second_0[43], y2[43], inv[0]);
    and s_143(second_1[43], y3[43], x[0]);
    and s_044(second_0[44], y2[44], inv[0]);
    and s_144(second_1[44], y3[44], x[0]);
    and s_045(second_0[45], y2[45], inv[0]);
    and s_145(second_1[45], y3[45], x[0]);
    and s_046(second_0[46], y2[46], inv[0]);
    and s_146(second_1[46], y3[46], x[0]);
    and s_047(second_0[47], y2[47], inv[0]);
    and s_147(second_1[47], y3[47], x[0]);
    and s_048(second_0[48], y2[48], inv[0]);
    and s_148(second_1[48], y3[48], x[0]);
    and s_049(second_0[49], y2[49], inv[0]);
    and s_149(second_1[49], y3[49], x[0]);
    and s_050(second_0[50], y2[50], inv[0]);
    and s_150(second_1[50], y3[50], x[0]);
    and s_051(second_0[51], y2[51], inv[0]);
    and s_151(second_1[51], y3[51], x[0]);
    and s_052(second_0[52], y2[52], inv[0]);
    and s_152(second_1[52], y3[52], x[0]);
    and s_053(second_0[53], y2[53], inv[0]);
    and s_153(second_1[53], y3[53], x[0]);
    and s_054(second_0[54], y2[54], inv[0]);
    and s_154(second_1[54], y3[54], x[0]);
    and s_055(second_0[55], y2[55], inv[0]);
    and s_155(second_1[55], y3[55], x[0]);
    and s_056(second_0[56], y2[56], inv[0]);
    and s_156(second_1[56], y3[56], x[0]);
    and s_057(second_0[57], y2[57], inv[0]);
    and s_157(second_1[57], y3[57], x[0]);
    and s_058(second_0[58], y2[58], inv[0]);
    and s_158(second_1[58], y3[58], x[0]);
    and s_059(second_0[59], y2[59], inv[0]);
    and s_159(second_1[59], y3[59], x[0]);
    and s_060(second_0[60], y2[60], inv[0]);
    and s_160(second_1[60], y3[60], x[0]);
    and s_061(second_0[61], y2[61], inv[0]);
    and s_161(second_1[61], y3[61], x[0]);
    and s_062(second_0[62], y2[62], inv[0]);
    and s_162(second_1[62], y3[62], x[0]);
    and s_063(second_0[63], y2[63], inv[0]);
    and s_163(second_1[63], y3[63], x[0]);

    wire[63 : 0] second;

    or s0(second[0], second_0[0], second_1[0]);
    or s1(second[1], second_0[1], second_1[1]);
    or s2(second[2], second_0[2], second_1[2]);
    or s3(second[3], second_0[3], second_1[3]);
    or s4(second[4], second_0[4], second_1[4]);
    or s5(second[5], second_0[5], second_1[5]);
    or s6(second[6], second_0[6], second_1[6]);
    or s7(second[7], second_0[7], second_1[7]);
    or s8(second[8], second_0[8], second_1[8]);
    or s9(second[9], second_0[9], second_1[9]);
    or s10(second[10], second_0[10], second_1[10]);
    or s11(second[11], second_0[11], second_1[11]);
    or s12(second[12], second_0[12], second_1[12]);
    or s13(second[13], second_0[13], second_1[13]);
    or s14(second[14], second_0[14], second_1[14]);
    or s15(second[15], second_0[15], second_1[15]);
    or s16(second[16], second_0[16], second_1[16]);
    or s17(second[17], second_0[17], second_1[17]);
    or s18(second[18], second_0[18], second_1[18]);
    or s19(second[19], second_0[19], second_1[19]);
    or s20(second[20], second_0[20], second_1[20]);
    or s21(second[21], second_0[21], second_1[21]);
    or s22(second[22], second_0[22], second_1[22]);
    or s23(second[23], second_0[23], second_1[23]);
    or s24(second[24], second_0[24], second_1[24]);
    or s25(second[25], second_0[25], second_1[25]);
    or s26(second[26], second_0[26], second_1[26]);
    or s27(second[27], second_0[27], second_1[27]);
    or s28(second[28], second_0[28], second_1[28]);
    or s29(second[29], second_0[29], second_1[29]);
    or s30(second[30], second_0[30], second_1[30]);
    or s31(second[31], second_0[31], second_1[31]);
    or s32(second[32], second_0[32], second_1[32]);
    or s33(second[33], second_0[33], second_1[33]);
    or s34(second[34], second_0[34], second_1[34]);
    or s35(second[35], second_0[35], second_1[35]);
    or s36(second[36], second_0[36], second_1[36]);
    or s37(second[37], second_0[37], second_1[37]);
    or s38(second[38], second_0[38], second_1[38]);
    or s39(second[39], second_0[39], second_1[39]);
    or s40(second[40], second_0[40], second_1[40]);
    or s41(second[41], second_0[41], second_1[41]);
    or s42(second[42], second_0[42], second_1[42]);
    or s43(second[43], second_0[43], second_1[43]);
    or s44(second[44], second_0[44], second_1[44]);
    or s45(second[45], second_0[45], second_1[45]);
    or s46(second[46], second_0[46], second_1[46]);
    or s47(second[47], second_0[47], second_1[47]);
    or s48(second[48], second_0[48], second_1[48]);
    or s49(second[49], second_0[49], second_1[49]);
    or s50(second[50], second_0[50], second_1[50]);
    or s51(second[51], second_0[51], second_1[51]);
    or s52(second[52], second_0[52], second_1[52]);
    or s53(second[53], second_0[53], second_1[53]);
    or s54(second[54], second_0[54], second_1[54]);
    or s55(second[55], second_0[55], second_1[55]);
    or s56(second[56], second_0[56], second_1[56]);
    or s57(second[57], second_0[57], second_1[57]);
    or s58(second[58], second_0[58], second_1[58]);
    or s59(second[59], second_0[59], second_1[59]);
    or s60(second[60], second_0[60], second_1[60]);
    or s61(second[61], second_0[61], second_1[61]);
    or s62(second[62], second_0[62], second_1[62]);
    or s63(second[63], second_0[63], second_1[63]);

    wire[63 : 0] result_0;
    wire[63 : 0] result_1;

    and r_00(result_0[0], first[0], inv[1]);
    and r_10(result_1[0], second[0], x[1]);
    and r_01(result_0[1], first[1], inv[1]);
    and r_11(result_1[1], second[1], x[1]);
    and r_02(result_0[2], first[2], inv[1]);
    and r_12(result_1[2], second[2], x[1]);
    and r_03(result_0[3], first[3], inv[1]);
    and r_13(result_1[3], second[3], x[1]);
    and r_04(result_0[4], first[4], inv[1]);
    and r_14(result_1[4], second[4], x[1]);
    and r_05(result_0[5], first[5], inv[1]);
    and r_15(result_1[5], second[5], x[1]);
    and r_06(result_0[6], first[6], inv[1]);
    and r_16(result_1[6], second[6], x[1]);
    and r_07(result_0[7], first[7], inv[1]);
    and r_17(result_1[7], second[7], x[1]);
    and r_08(result_0[8], first[8], inv[1]);
    and r_18(result_1[8], second[8], x[1]);
    and r_09(result_0[9], first[9], inv[1]);
    and r_19(result_1[9], second[9], x[1]);
    and r_010(result_0[10], first[10], inv[1]);
    and r_110(result_1[10], second[10], x[1]);
    and r_011(result_0[11], first[11], inv[1]);
    and r_111(result_1[11], second[11], x[1]);
    and r_012(result_0[12], first[12], inv[1]);
    and r_112(result_1[12], second[12], x[1]);
    and r_013(result_0[13], first[13], inv[1]);
    and r_113(result_1[13], second[13], x[1]);
    and r_014(result_0[14], first[14], inv[1]);
    and r_114(result_1[14], second[14], x[1]);
    and r_015(result_0[15], first[15], inv[1]);
    and r_115(result_1[15], second[15], x[1]);
    and r_016(result_0[16], first[16], inv[1]);
    and r_116(result_1[16], second[16], x[1]);
    and r_017(result_0[17], first[17], inv[1]);
    and r_117(result_1[17], second[17], x[1]);
    and r_018(result_0[18], first[18], inv[1]);
    and r_118(result_1[18], second[18], x[1]);
    and r_019(result_0[19], first[19], inv[1]);
    and r_119(result_1[19], second[19], x[1]);
    and r_020(result_0[20], first[20], inv[1]);
    and r_120(result_1[20], second[20], x[1]);
    and r_021(result_0[21], first[21], inv[1]);
    and r_121(result_1[21], second[21], x[1]);
    and r_022(result_0[22], first[22], inv[1]);
    and r_122(result_1[22], second[22], x[1]);
    and r_023(result_0[23], first[23], inv[1]);
    and r_123(result_1[23], second[23], x[1]);
    and r_024(result_0[24], first[24], inv[1]);
    and r_124(result_1[24], second[24], x[1]);
    and r_025(result_0[25], first[25], inv[1]);
    and r_125(result_1[25], second[25], x[1]);
    and r_026(result_0[26], first[26], inv[1]);
    and r_126(result_1[26], second[26], x[1]);
    and r_027(result_0[27], first[27], inv[1]);
    and r_127(result_1[27], second[27], x[1]);
    and r_028(result_0[28], first[28], inv[1]);
    and r_128(result_1[28], second[28], x[1]);
    and r_029(result_0[29], first[29], inv[1]);
    and r_129(result_1[29], second[29], x[1]);
    and r_030(result_0[30], first[30], inv[1]);
    and r_130(result_1[30], second[30], x[1]);
    and r_031(result_0[31], first[31], inv[1]);
    and r_131(result_1[31], second[31], x[1]);
    and r_032(result_0[32], first[32], inv[1]);
    and r_132(result_1[32], second[32], x[1]);
    and r_033(result_0[33], first[33], inv[1]);
    and r_133(result_1[33], second[33], x[1]);
    and r_034(result_0[34], first[34], inv[1]);
    and r_134(result_1[34], second[34], x[1]);
    and r_035(result_0[35], first[35], inv[1]);
    and r_135(result_1[35], second[35], x[1]);
    and r_036(result_0[36], first[36], inv[1]);
    and r_136(result_1[36], second[36], x[1]);
    and r_037(result_0[37], first[37], inv[1]);
    and r_137(result_1[37], second[37], x[1]);
    and r_038(result_0[38], first[38], inv[1]);
    and r_138(result_1[38], second[38], x[1]);
    and r_039(result_0[39], first[39], inv[1]);
    and r_139(result_1[39], second[39], x[1]);
    and r_040(result_0[40], first[40], inv[1]);
    and r_140(result_1[40], second[40], x[1]);
    and r_041(result_0[41], first[41], inv[1]);
    and r_141(result_1[41], second[41], x[1]);
    and r_042(result_0[42], first[42], inv[1]);
    and r_142(result_1[42], second[42], x[1]);
    and r_043(result_0[43], first[43], inv[1]);
    and r_143(result_1[43], second[43], x[1]);
    and r_044(result_0[44], first[44], inv[1]);
    and r_144(result_1[44], second[44], x[1]);
    and r_045(result_0[45], first[45], inv[1]);
    and r_145(result_1[45], second[45], x[1]);
    and r_046(result_0[46], first[46], inv[1]);
    and r_146(result_1[46], second[46], x[1]);
    and r_047(result_0[47], first[47], inv[1]);
    and r_147(result_1[47], second[47], x[1]);
    and r_048(result_0[48], first[48], inv[1]);
    and r_148(result_1[48], second[48], x[1]);
    and r_049(result_0[49], first[49], inv[1]);
    and r_149(result_1[49], second[49], x[1]);
    and r_050(result_0[50], first[50], inv[1]);
    and r_150(result_1[50], second[50], x[1]);
    and r_051(result_0[51], first[51], inv[1]);
    and r_151(result_1[51], second[51], x[1]);
    and r_052(result_0[52], first[52], inv[1]);
    and r_152(result_1[52], second[52], x[1]);
    and r_053(result_0[53], first[53], inv[1]);
    and r_153(result_1[53], second[53], x[1]);
    and r_054(result_0[54], first[54], inv[1]);
    and r_154(result_1[54], second[54], x[1]);
    and r_055(result_0[55], first[55], inv[1]);
    and r_155(result_1[55], second[55], x[1]);
    and r_056(result_0[56], first[56], inv[1]);
    and r_156(result_1[56], second[56], x[1]);
    and r_057(result_0[57], first[57], inv[1]);
    and r_157(result_1[57], second[57], x[1]);
    and r_058(result_0[58], first[58], inv[1]);
    and r_158(result_1[58], second[58], x[1]);
    and r_059(result_0[59], first[59], inv[1]);
    and r_159(result_1[59], second[59], x[1]);
    and r_060(result_0[60], first[60], inv[1]);
    and r_160(result_1[60], second[60], x[1]);
    and r_061(result_0[61], first[61], inv[1]);
    and r_161(result_1[61], second[61], x[1]);
    and r_062(result_0[62], first[62], inv[1]);
    and r_162(result_1[62], second[62], x[1]);
    and r_063(result_0[63], first[63], inv[1]);
    and r_163(result_1[63], second[63], x[1]);

    or r0(z[0], result_0[0], result_1[0]);
    or r1(z[1], result_0[1], result_1[1]);
    or r2(z[2], result_0[2], result_1[2]);
    or r3(z[3], result_0[3], result_1[3]);
    or r4(z[4], result_0[4], result_1[4]);
    or r5(z[5], result_0[5], result_1[5]);
    or r6(z[6], result_0[6], result_1[6]);
    or r7(z[7], result_0[7], result_1[7]);
    or r8(z[8], result_0[8], result_1[8]);
    or r9(z[9], result_0[9], result_1[9]);
    or r10(z[10], result_0[10], result_1[10]);
    or r11(z[11], result_0[11], result_1[11]);
    or r12(z[12], result_0[12], result_1[12]);
    or r13(z[13], result_0[13], result_1[13]);
    or r14(z[14], result_0[14], result_1[14]);
    or r15(z[15], result_0[15], result_1[15]);
    or r16(z[16], result_0[16], result_1[16]);
    or r17(z[17], result_0[17], result_1[17]);
    or r18(z[18], result_0[18], result_1[18]);
    or r19(z[19], result_0[19], result_1[19]);
    or r20(z[20], result_0[20], result_1[20]);
    or r21(z[21], result_0[21], result_1[21]);
    or r22(z[22], result_0[22], result_1[22]);
    or r23(z[23], result_0[23], result_1[23]);
    or r24(z[24], result_0[24], result_1[24]);
    or r25(z[25], result_0[25], result_1[25]);
    or r26(z[26], result_0[26], result_1[26]);
    or r27(z[27], result_0[27], result_1[27]);
    or r28(z[28], result_0[28], result_1[28]);
    or r29(z[29], result_0[29], result_1[29]);
    or r30(z[30], result_0[30], result_1[30]);
    or r31(z[31], result_0[31], result_1[31]);
    or r32(z[32], result_0[32], result_1[32]);
    or r33(z[33], result_0[33], result_1[33]);
    or r34(z[34], result_0[34], result_1[34]);
    or r35(z[35], result_0[35], result_1[35]);
    or r36(z[36], result_0[36], result_1[36]);
    or r37(z[37], result_0[37], result_1[37]);
    or r38(z[38], result_0[38], result_1[38]);
    or r39(z[39], result_0[39], result_1[39]);
    or r40(z[40], result_0[40], result_1[40]);
    or r41(z[41], result_0[41], result_1[41]);
    or r42(z[42], result_0[42], result_1[42]);
    or r43(z[43], result_0[43], result_1[43]);
    or r44(z[44], result_0[44], result_1[44]);
    or r45(z[45], result_0[45], result_1[45]);
    or r46(z[46], result_0[46], result_1[46]);
    or r47(z[47], result_0[47], result_1[47]);
    or r48(z[48], result_0[48], result_1[48]);
    or r49(z[49], result_0[49], result_1[49]);
    or r50(z[50], result_0[50], result_1[50]);
    or r51(z[51], result_0[51], result_1[51]);
    or r52(z[52], result_0[52], result_1[52]);
    or r53(z[53], result_0[53], result_1[53]);
    or r54(z[54], result_0[54], result_1[54]);
    or r55(z[55], result_0[55], result_1[55]);
    or r56(z[56], result_0[56], result_1[56]);
    or r57(z[57], result_0[57], result_1[57]);
    or r58(z[58], result_0[58], result_1[58]);
    or r59(z[59], result_0[59], result_1[59]);
    or r60(z[60], result_0[60], result_1[60]);
    or r61(z[61], result_0[61], result_1[61]);
    or r62(z[62], result_0[62], result_1[62]);
    or r63(z[63], result_0[63], result_1[63]);

endmodule
